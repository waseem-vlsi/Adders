
module adder(
input a,b,c,
output p,g,s);
 
 assign g = a&b;
 assign p = a^b;
 assign s = a^b^c; 
endmodule
module carry_gen(
input [3:0]p,g,
input cin,
output cout,P0,G0,
output c1,c2,c3,c4);
wire c4;
assign c1 = g[0]|(p[0]&cin), c2 = g[1]|(p[1]&g[0])|(p[1]&p[0]&cin) , c3 = g[2]| (p[2]&g[1])|(p[2]&p[1]&g[0])|(p[2]&p[1]&p[0]&cin),  c4 = g[3]|(p[3]&g[2])| (p[3]&g[2]&g[1])|(p[3]&p[2]&p[1]&g[0])|(p[3]&p[2]&p[1]&p[0]&cin);
assign P0 = p[3] & p[2] & p[1] & p[0], G0 = g[3] | (p[3] &g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]); 
assign cout = c4;
endmodule

module  CLA_4_bit(
input [3:0]a,b,
input cin,
output [3:0]sum,
output cout);
wire [3:0]p,g;
wire c1,c2,c3,c4,P0,G0;
adder A1(.a(a[0]), .b(b[0]), .s(sum[0]),.p(p[0]), .g(g[0]), .c(cin));
adder A2(.a(a[1]), .b(b[1]), .s(sum[1]),.p(p[1]), .g(g[1]), .c(c1));
adder A3(.a(a[2]), .b(b[2]), .s(sum[2]),.p(p[2]), .g(g[2]), .c(c2));
adder A4(.a(a[3]), .b(b[3]), .s(sum[3]),.p(p[3]), .g(g[3]),.c(c3));
carry_gen A5(.p(p), .g(g), .c1(c1), .c2(c2),.c3(c3), .c4(cout), .P0(P0), .G0(G0), .cin(cin));
endmodule


// MAIN MODULE


module hybrid_RCA_CLA_12_bit(
input [11:0]A,B,
input Cin,
output [12:0]Y);
wire carry1,carry2;
wire [11:0]S;
wire carry,C;
 CLA_4_bit A1(.a(A[3:0]), .b(B[3:0]), .cin(Cin), .sum(S[3:0]), .cout(carry1));
 CLA_4_bit A2(.a(A[7:4]), .b(B[7:4]), .cin(carry1), .sum(S[7:4]), .cout(carry2));
 CLA_4_bit A3(.a(A[11:8]), .b(B[11:8]), .cin(carry2), .sum(S[11:8]), .cout(C));
 assign Y = {C,S}; 
endmodule
