`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

module RCA_4bit_tb( );
reg [3:0]a,b;
reg cin;
wire [3:0]sum;
wire cout;
RCA_4bit DUT(.a(a), .b(b), .cin(cin), .sum(sum), .cout(cout));
initial
begin
#10 a = 4'b0000; b = 4'b0001; cin = 4'b0000;
#10 a = 4'b0001; b = 4'b0001; cin = 4'b0000;
#10 a = 4'b0000; b = 4'b0001; cin = 4'b0000;
#10 a = 4'b0001; b = 4'b0001; cin = 4'b0101;
#10 a = 4'b1111; b = 4'b0111; cin = 4'b0010;
#5 $finish;
end
endmodule

