`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////


module RCA_16bit_tb();
reg [15:0]a,b;
reg cin;
wire [15:0]sum;
wire cout;
RCA_16bit DUT(.a(a), .b(b), .cin(cin), .sum(sum), .cout(cout));
initial
begin
#10 cin = 1'b0;
#10 a = 16'b0000000000000000; b = 4'b0000000000001111; 
#10 a = 16'b0000000000000010; b = 4'b0000000000001110; 
#10 a = 16'b0000000000000010; b = 4'b0000000000000011; 
#10 a = 16'b0000000000000001; b = 4'b0000000000001111; 
#10 a = 16'b0000000000000001; b = 4'b0000000000000011;
#10 a = 16'b0000000000000000; b = 4'b0000000000001111; 

#5 $finish;
end
endmodule
